package synch_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "sequence_item.svh"
    `include "random_sequence.svh"    
    `include "write_sequence.svh"
    `include "read_sequence.svh"    
    `include "sequencer.svh"
    `include "driver.svh"    
    `include "monitor.svh"   
    `include "agent.svh"   
    `include "scoreboard.svh"   
    `include "coverage.svh"     
    `include "env.svh"   
    `include "SerialSeq.svh"
    `include "full_test.svh" 
endpackage :synch_pkg