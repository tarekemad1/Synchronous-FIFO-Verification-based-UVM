package SynchFifo_pkg;
    import uvm_pkg ::*;
    import SynchFifo_pkg::*;
    `include "uvm_macros.svh";
    `include "sequence_item.svh";
    `include "sequencer.svh";
    `include "base_sequence.svh";
    `include "monitor.svh";
    `include "agent.svh";
    `include "coverage.svh";
    `include "env.svh";
    `include "base_test.svh";
    
    
endpackage